library verilog;
use verilog.vl_types.all;
entity sdram_controller_tb is
end sdram_controller_tb;
