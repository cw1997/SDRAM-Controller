library verilog;
use verilog.vl_types.all;
entity auto_refresh_counter_tb is
end auto_refresh_counter_tb;
